
library IEEE;
use IEEE.std_logic_1164.all;


package array_package_0to1 is
	type vector_array_0to1 is array (0 to 0) of std_logic_vector(31 downto 0);
end package array_package_0to1;
library IEEE;
use IEEE.std_logic_1164.all;


package mux2to1_array_package is
	type size2_vector_array is array (0 to 1) of std_logic_vector(31 downto 0);
end package mux2to1_array_package;


library IEEE;
use IEEE.std_logic_1164.all;

entity dec5to32 is
	
	port(i_S : in std_logic_vector(4 downto 0);
	     i_EN : std_logic;
	     o_Q : out std_logic_vector(31 downto 0));

end dec5to32;

architecture dataflow of dec5to32 is

begin

    process(i_S, i_EN)
    begin
        if i_EN = '1' then
            case i_S is
                when "00000" => o_Q <= "00000000000000000000000000000001";
                when "00001" => o_Q <= "00000000000000000000000000000010";
                when "00010" => o_Q <= "00000000000000000000000000000100";
                when "00011" => o_Q <= "00000000000000000000000000001000";
                when "00100" => o_Q <= "00000000000000000000000000010000";
                when "00101" => o_Q <= "00000000000000000000000000100000";
                when "00110" => o_Q <= "00000000000000000000000001000000";
                when "00111" => o_Q <= "00000000000000000000000010000000";
                when "01000" => o_Q <= "00000000000000000000000100000000";
                when "01001" => o_Q <= "00000000000000000000001000000000";
                when "01010" => o_Q <= "00000000000000000000010000000000";
                when "01011" => o_Q <= "00000000000000000000100000000000";
                when "01100" => o_Q <= "00000000000000000001000000000000";
                when "01101" => o_Q <= "00000000000000000010000000000000";
                when "01110" => o_Q <= "00000000000000000100000000000000";
                when "01111" => o_Q <= "00000000000000001000000000000000";
                when "10000" => o_Q <= "00000000000000010000000000000000";
                when "10001" => o_Q <= "00000000000000100000000000000000";
                when "10010" => o_Q <= "00000000000001000000000000000000";
                when "10011" => o_Q <= "00000000000010000000000000000000";
                when "10100" => o_Q <= "00000000000100000000000000000000";
                when "10101" => o_Q <= "00000000001000000000000000000000";
                when "10110" => o_Q <= "00000000010000000000000000000000";
                when "10111" => o_Q <= "00000000100000000000000000000000";
                when "11000" => o_Q <= "00000001000000000000000000000000";
                when "11001" => o_Q <= "00000010000000000000000000000000";
                when "11010" => o_Q <= "00000100000000000000000000000000";
                when "11011" => o_Q <= "00001000000000000000000000000000";
                when "11100" => o_Q <= "00010000000000000000000000000000";
                when "11101" => o_Q <= "00100000000000000000000000000000";
                when "11110" => o_Q <= "01000000000000000000000000000000";
                when "11111" => o_Q <= "10000000000000000000000000000000";
                when others  => o_Q <= "00000000000000000000000000000000"; --debug
            end case;
        else
            o_Q <= "00000000000000000000000000000000"; -- disabled
        end if;
    end process;

end dataflow;

